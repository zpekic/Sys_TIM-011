----------------------------------------------------------------------------------
-- Company: @Home
-- Engineer: zpekic@hotmail.com
-- 
-- Create Date: 08/29/2020 11:13:02 PM
-- Design Name: Various TIM-011 components
-- Module Name: sys_tim-011_mercury - Behavioral
-- Project Name: 
-- Target Devices: https://www.micro-nova.com/mercury/ + Baseboard
-- Input devices: 
--
-- Tool Versions: ISE 14.7 (nt)
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.99 - Kinda works...
-- Additional Comments:
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
--use work.tms0800_package.all;

entity sys_tim011_mercury is
    Port ( 
				-- 50MHz on the Mercury board
				CLK: in std_logic;
				
				-- 12MHz external clock
				EXT_CLK: in std_logic;
				
				-- Master reset button on Mercury board
				USR_BTN: in std_logic; 

				-- Switches on baseboard
				-- SW(0) -- direction when scrolling
				-- SW(1) -- data source selection for 7seg display
				-- SW(2) -- palette selection (best on)
				-- SW(3) -- palette selection (best off)
				-- SW(4) -- off
				-- SW(5) -- on
				-- SW(6) -- off
				-- SW(7)	-- off

				SW: in std_logic_vector(7 downto 0); 

				-- Push buttons on baseboard
				-- BTN0 - scroll
				-- BTN1 - video only test pattern (memory not affected)
				-- BTN2 - fill left/right
				-- BTN3 - fill top/down
				BTN: in std_logic_vector(3 downto 0); 

				-- Stereo audio output on baseboard
				AUDIO_OUT_L, AUDIO_OUT_R: out std_logic;

				-- 7seg LED on baseboard 
				A_TO_G: out std_logic_vector(6 downto 0); 
				AN: out std_logic_vector(3 downto 0); 
				DOT: out std_logic; 
				-- 4 LEDs on Mercury board (3 and 2 are used by VGA VSYNC and HSYNC)
				LED: inout std_logic_vector(3 downto 0);

				-- ADC interface
				-- channel	input
				-- 0			Audio Left
				-- 1 			Audio Right
				-- 2			Temperature
				-- 3			Light	
				-- 4			Pot
				-- 5			Channel 5 (free)
				-- 6			Channel 6 (free)
				-- 7			Channel 7 (free)
				ADC_MISO: in std_logic;
				ADC_MOSI: out std_logic;
				ADC_SCK: out std_logic;
				ADC_CSN: out std_logic;
				--PS2_DATA: in std_logic;
				--PS2_CLOCK: in std_logic;

				--VGA interface
				--register state is traced to VGA after each instruction if SW0 = on
				--640*480 50Hz mode is used, which give 80*60 character display
				--but to save memory, only 80*50 are used which fits into 4k video RAM
				--HSYNC: out std_logic;
				--VSYNC: out std_logic;
				--RED: out std_logic_vector(2 downto 0);
				--GRN: out std_logic_vector(2 downto 0);
				--BLU: out std_logic_vector(1 downto 0);
				
				--PMOD interface
				--connection to https://store.digilentinc.com/pmod-kypd-16-button-keypad/
				PMOD: inout std_logic_vector(7 downto 0)
          );
end sys_tim011_mercury;

architecture Structural of sys_tim011_mercury is

component Grafika is
    Port ( -- 
	 		  dotclk : in  STD_LOGIC;
           a : in  STD_LOGIC_VECTOR (15 downto 0);
           nRD : in  STD_LOGIC;
           nWR : in  STD_LOGIC;
           d : inout  STD_LOGIC_VECTOR (7 downto 0);
           ioe : in  STD_LOGIC;
           nScroll : in  STD_LOGIC;
			  -- debug
			  test: in STD_LOGIC;
			  vid_gated: STD_LOGIC;
			  -- monitor side
			  hsync: out STD_LOGIC;
			  vsync: out STD_LOGIC;
			  vid1: out STD_LOGIC;
			  vid2: out STD_LOGIC
			);
end component;

component oneshot is
    Port ( trigger : in  STD_LOGIC;
           tick : in  STD_LOGIC;
           duration : in  STD_LOGIC_VECTOR (15 downto 0);
           shot : out  STD_LOGIC);
end component;

component sn74ls283 is
    Port ( c0 : in  STD_LOGIC;
           a : in  STD_LOGIC_VECTOR (4 downto 1);
           b : in  STD_LOGIC_VECTOR (4 downto 1);
           s : out  STD_LOGIC_VECTOR (4 downto 1);
           c4 : out  STD_LOGIC);
end component;

component sn74ls374 is
    Port ( nOC : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           D : in  STD_LOGIC_VECTOR (7 downto 0);
           Q : out  STD_LOGIC_VECTOR (7 downto 0));
end component;

component sn74hc4040 is
    Port ( q12_1 : out  STD_LOGIC;
           q6_2 : out  STD_LOGIC;
           q5_3 : out  STD_LOGIC;
           q7_4 : out  STD_LOGIC;
           q4_5 : out  STD_LOGIC;
           q3_6 : out  STD_LOGIC;
           q2_7 : out  STD_LOGIC;
           q1_9 : out  STD_LOGIC;
           clock_10 : in  STD_LOGIC;
           reset_11 : in  STD_LOGIC;
           q9_12 : out  STD_LOGIC;
           q8_13 : out  STD_LOGIC;
           q10_14 : out  STD_LOGIC;
           q11_15 : out  STD_LOGIC);
end component;

component fourdigitsevensegled is
    Port ( -- inputs
			  hexdata : in  STD_LOGIC_VECTOR (3 downto 0);
           digsel : in  STD_LOGIC_VECTOR (1 downto 0);
           showdigit : in  STD_LOGIC_VECTOR (3 downto 0);
           showdot : in  STD_LOGIC_VECTOR (3 downto 0);
			  -- outputs
           anode : out  STD_LOGIC_VECTOR (3 downto 0);
           segment : out  STD_LOGIC_VECTOR (7 downto 0)
			 );
end component;

component interactivereg is
    Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           enable : in  STD_LOGIC;
           init : in  STD_LOGIC_VECTOR (15 downto 0);
           up : in  STD_LOGIC;
           down : in  STD_LOGIC;
           value : buffer  STD_LOGIC_VECTOR (15 downto 0));
end component;

--component mouse_ctrl is
--  generic (
--    X_MAX : integer := 799; -- maximum X position
--    Y_MAX : integer := 599  -- maximum Y position
--    );
--  port(
--    clk25        : in    std_logic;                 -- 25MHz clock
--    clr          : in    std_logic;                 -- async clear
--    PS2C         : inout std_logic;                 -- PS/2 clock
--    PS2D         : inout std_logic;                 -- PS/2 data
--    click_middle : out   std_logic;                 -- middle click
--    click_right  : out   std_logic;                 -- right click
--    click_left   : out   std_logic;                 -- left click
--    x_position   : out   integer range 0 to X_MAX;  -- current X position
--    y_position   : out   integer range 0 to Y_MAX   -- current Y position
--    );
--end component;

component freqcounter is
    Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           freq : in  STD_LOGIC;
			  bcd:	in STD_LOGIC;
           value : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component uart_receiver is
    Port ( rx_clk4 : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           rx : in  STD_LOGIC;
           mode : in  STD_LOGIC_VECTOR (2 downto 0);
			  frame_active: out  STD_LOGIC;
           frame_ready : out  STD_LOGIC;
           frame_valid : out  STD_LOGIC;
           frame_data : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component signalcounter is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           input : in  STD_LOGIC;
           sel : in  STD_LOGIC;
           count : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component configurabledelayline is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           init : in  STD_LOGIC;
           delay : in  STD_LOGIC_VECTOR (3 downto 0);
           signal_in : in  STD_LOGIC;
           signal_out : out  STD_LOGIC);
end component;

--component rx_reg is
--    Port ( clk : in  STD_LOGIC;
--           reset : in  STD_LOGIC;
--           enable : in  STD_LOGIC;
--           rx : in  STD_LOGIC;
--           d : out  STD_LOGIC_VECTOR (7 downto 0);
--           dready : out  STD_LOGIC);
--end component;

component ps2tim is
    Port ( reset : in  STD_LOGIC;
           uart_clk4 : in  STD_LOGIC;
           uart_rx : in  STD_LOGIC;
           uart_tx : out  STD_LOGIC;
           ps2_clk : inout  STD_LOGIC;
           ps2_data : inout  STD_LOGIC;
			  debugsel: in STD_LOGIC;
           debug : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component debouncer8channel is
    Port ( clock : in STD_LOGIC;
           reset : in STD_LOGIC;
           signal_raw : in STD_LOGIC_VECTOR (7 downto 0);
           signal_debounced : out STD_LOGIC_VECTOR (7 downto 0));
end component;

component memconsole is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           control : in  STD_LOGIC_VECTOR (3 downto 0);
           EN : out  STD_LOGIC;
           RD : out  STD_LOGIC;
           WR : out  STD_LOGIC;
           A : out  STD_LOGIC_VECTOR (15 downto 0);
           D : inout  STD_LOGIC_VECTOR (7 downto 0);
           DD : out  STD_LOGIC_VECTOR (7 downto 0));
end component;

component memtester is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
			  fill: in STD_LOGIC;
			  direction: in STD_LOGIC;
           EN : out  STD_LOGIC;
           RD : out  STD_LOGIC;
           WR : out  STD_LOGIC;
           A : out  STD_LOGIC_VECTOR (15 downto 0);
           D : inout  STD_LOGIC_VECTOR (7 downto 0);
           DD : out  STD_LOGIC_VECTOR (7 downto 0));
end component;

type palette is array (0 to 15) of std_logic_vector(2 downto 0);
signal bgr: palette := (
	"011",	-- yellow -- this palette looks bad probably because base background color is not black
	"110",	-- cyan
	"101",	-- purple
	"111",	-- white

	"000",	-- black
	"101",	-- purple
	"110",	-- cyan
	"100",	-- blue

	"000",	-- black
	"011",	-- yellow
	"110",	-- cyan
	"010",	-- green

	"000",	-- black
	"011",	-- yellow
	"101",	-- purple
	"001" 	-- red
);

signal RESET: std_logic;

-- debug
signal test_static, test_dynamic, test_scroll, test_clk, nScrollEnable: std_logic;
signal digsel: std_logic_vector(1 downto 0);
signal offset_new: std_logic_vector(7 downto 0);
signal offset_add_lo_cout: std_logic;
--signal h, digsel0_delayed: std_logic;
signal hexdata, hexsel, showdigit: std_logic_vector(3 downto 0);
---
signal data: std_logic_vector(15 downto 0);
signal freq_uart, freq_uart4: std_logic;

--- frequency signals
signal freq24M, dotclk: std_logic;
signal prescale_baud, prescale_power: integer range 0 to 65535;
signal freq153600, freq76800, freq38400, freq19200, freq9600, freq4800, freq2400, freq1200, freq600, freq300: std_logic;		
signal freq4096, freq2, freq4: std_logic;		

--- video sync signals
signal gr_hsync, gr_vsync: std_logic;
signal sh_hsync, sh_vsync : std_logic;
signal out_hsync, out_vsync : std_logic;
signal hsync_cnt, vsync_cnt, h_duration, v_duration: std_logic_vector(15 downto 0); 
signal enable_hshot, enable_vshot : std_logic;
-- video data signals
signal gr_vid2, gr_vid1: std_logic;
signal color: std_logic_vector(3 downto 0); -- combines one of 1 palettes plus vid2 and vid1
-- video memory bus
signal vm_en, vm_rd, vm_wr: std_logic;
signal D, DD: std_logic_vector(7 downto 0);
signal A: std_logic_vector(15 downto 0);

---
signal switch, button: std_logic_vector(7 downto 0);
--- test mouse
--signal mouse_left, mouse_right, mouse_middle: std_logic;
--signal mouse_x: integer range 0 to 511;
--signal mouse_y: integer range 0 to 255;

--alias ps2_data: std_logic is LED(0);
--alias ps2_clk: std_logic is LED(1);
--signal frame_parity: std_logic;

-- ADC
signal adc_trigger  : std_logic := '1';              -- go sample from ADC
signal adc_done     : std_logic := '0';              -- done sampling ADC
signal adc_dout     : std_logic_vector(9 downto 0);  -- ADC data out
signal adc_data_reg : unsigned(9 downto 0);          -- ADC data registered
signal adc_channel  : std_logic_vector(2 downto 0);  -- ADC channel
signal adc_clk: std_logic;
signal min: unsigned(9 downto 0) := "1111111111";
signal max: unsigned(9 downto 0) := "0000000000";
signal adc_count, adc_old_count, freq_value: std_logic_vector(15 downto 0);
signal adc_value: std_logic_vector(7 downto 0);
signal f_in, f_out, f_in_audio: std_logic;
-- UART
signal frame_ready, frame_valid, frame_active: std_logic;
signal frame_data, uart_frame, display: std_logic_vector(15 downto 0);
signal rx, rx_analog, rx_digital: std_logic;
signal baudrate_x1, baudrate_x2, baudrate_x4: std_logic;
signal sr: std_logic_vector(31 downto 0);
  
begin
   
RESET <= USR_BTN;
--dotclk <= EXT_CLK;	-- 12MHz "half-size" crystal on Mercury baseboard
	
clockgen: sn74hc4040 port map (
			clock_10 => EXT_CLK,	-- 48MHz "half-size" crystal on Mercury baseboard
			reset_11 => RESET,
			q1_9 => freq24M, 
			q2_7 => dotclk,
			q3_6 => open, --PMOD(7),		-- 6.25
			q4_5 => open, --PMOD(6),		-- 3.125
			q5_3 => open, --PMOD(5),		-- 1.5625
			q6_2 => open, --PMOD(4), 		-- 0.78125
			q7_4 =>   open,		-- 0.390625
			q8_13 =>  open,		-- 0.1953125
			q9_12 =>  open,		-- 0.09765625
			q10_14 => open,		-- 0.048828125
			q11_15 => digsel(0),	-- 0.0244140625
			q12_1 =>  digsel(1)	-- 0.01220703125
		);
--
prescale: process(CLK, freq153600, freq4096)
begin
	if (rising_edge(CLK)) then
		if (prescale_baud = 0) then
			freq153600 <= not freq153600;
			prescale_baud <= (50000000 / (2 * 153600));
		else
			prescale_baud <= prescale_baud - 1;
		end if;
		if (prescale_power = 0) then
			freq4096 <= not freq4096;
			prescale_power <= (50000000 / (2 * 4096));
		else
			prescale_power <= prescale_power - 1;
		end if;
	end if;
end process;
--
baudgen: sn74hc4040 port map (
			clock_10 => freq153600,
			reset_11 => RESET,
			q1_9 => freq76800, 
			q2_7 => freq38400,
			q3_6 => freq19200,		
			q4_5 => freq9600,		
			q5_3 => freq4800,		
			q6_2 => freq2400, 	
			q7_4 => freq1200,		
			q8_13 => freq600,		
			q9_12 =>  freq300,
			q10_14 => open,	
			q11_15 => open,	
			q12_1 =>  open	
		);
--
powergen: sn74hc4040 port map (
			clock_10 => freq4096,
			reset_11 => RESET,
			q1_9 => open, 
			q2_7 => open,
			q3_6 => open,		
			q4_5 => open,		
			q5_3 => open,		
			q6_2 => open, 	
			q7_4 => open,		
			q8_13 => open,		
			q9_12 =>  open,	
			q10_14 => freq4,	
			q11_15 => freq2,	
			q12_1 =>  open	
		);
--	
	debounce_sw: debouncer8channel Port map ( 
		clock => freq19200, 
		reset => RESET,
		signal_raw => SW,
		signal_debounced => switch
	);

	debounce_btn: debouncer8channel Port map ( 
		clock => freq19200, 
		reset => RESET,
		signal_raw(7 downto 4) => "0000",
		signal_raw(3 downto 0) => BTN,
		signal_debounced => button
	);
	
kbd: ps2tim Port map ( 
			reset => RESET,
         uart_clk4 => freq38400, -- baudrate = /4 = 9600
         uart_rx => '1', --PMOD(5),		-- TODO: verify pin
         uart_tx => open, --PMOD(6),		-- TODO: verify pin
         ps2_clk => LED(1),
         ps2_data => LED(0),
			debugsel => switch(0),
         debug => open--display
		);
	
--  -- mouse controller
--  mouse : entity work.mouse_ctrl
--    generic map (
--      X_MAX => 511,
--      Y_MAX => 255
--      )
--    port map(
--      clk25        => freq25M,
--      clr          => '0',
--      PS2C         => ps2_clk,
--      PS2D         => ps2_data,
--      click_middle => mouse_middle,
--      click_right  => mouse_right,
--      click_left   => mouse_left,
--      x_position   => mouse_x,
--      y_position   => mouse_y
--      );
--		
--console: memconsole Port map(
--			clk => freq2,
--         reset => RESET,
--         control => button(3 downto 0),
--         EN => vm_en,
--         RD => vm_rd,
--         WR => vm_wr,
--         A => A,
--         D => D,
--         DD => DD
--	);

mtest: memtester Port map(
			clk => test_clk,
         reset => RESET,
			fill => test_dynamic,
			direction => button(2),
         EN => vm_en,
         RD => vm_rd,
         WR => vm_wr,
         A => A,
         D => D,
         DD => DD
	);
--	
test_static <= '1' when (button(3 downto 0) = "0010") else '0';
test_dynamic <= '0' when (button(3 downto 2) = "00") else '1';
test_scroll <= nScrollEnable when (button(3 downto 0) = "0001") else '1';

test_clk <= freq38400 when (button(3 downto 2) = "11") else freq9600;

-- scroll logic
nScrollEnable <= vm_en or vm_rd or vm_wr;	-- low if all all, meaning no other bus activity

offset_reg: sn74ls374 Port map ( 
			nOC => nScrollEnable,
         CLK => test_scroll,
         D => offset_new,
         Q => D
	);

offset_add_hi: sn74ls283 Port map ( -- add +1 or -1 to offset)
			c0 => offset_add_lo_cout,
			a(4) => switch(0),
			a(3) => switch(0),
			a(2) => switch(0),
			a(1) => switch(0),
			b => D(7 downto 4),
			s => offset_new(7 downto 4),
			c4 => open
	);
	
offset_add_lo: sn74ls283 Port map ( 
			c0 => '0',
			a(4) => switch(0),
			a(3) => switch(0),
			a(2) => switch(0),
			a(1) => '1',
			b => D(3 downto 0),
			s => offset_new(3 downto 0),
			c4 => offset_add_lo_cout
	);	
--	

	video: Grafika port map (
		-- system
		  dotclk => dotclk,
		  A(15) => '1',	-- mapped to 0x8000 - 0xFFFF or extended IO space
		  A(14 downto 0) => A(14 downto 0),
		  nRD => not (vm_rd),
		  nWR => not (vm_wr),
		  d => D,
		  ioe => vm_en,
		  nScroll => test_scroll,
		-- debug
		  test => test_static,
		  vid_gated => '0', -- do not gate vid1/2 on dotclk (this is different from original!)
		-- monitor side
		  hsync => gr_hsync, --HSYNC,
		  vsync => gr_vsync,--VSYNC,
		  vid1 => gr_vid1, --BLU(0),
		  vid2 => gr_vid2  --BLU(1)
	);
	
--LED(0) <= dotclk;
--LED(1) <= vm_en;
LED(2) <= vm_rd;
LED(3) <= vm_wr;

-- Connect to GBS8200 gray wire
	PMOD(3) <= out_hsync xor out_vsync;
	
-- connect to GBS8200 blue / green / red wires
	PMOD(2 downto 0) <= bgr(to_integer(unsigned(color)));
	color <= switch(3 downto 2) & gr_vid2 & gr_vid1;

--	HSYNC <= not sh_hsync;
--	VSYNC <= not sh_vsync;
--	BLU(1) <= switch(1) xor gr_vid2;
--	BLU(0) <= switch(0) xor gr_vid1;
--	RED <= "000";
--	GRN <= "000";

--with switch(7 downto 6) select
		out_hsync <= 	gr_hsync; -- when "00",
							--sh_hsync when "01",
							--not gr_hsync when "10",			-- STABLE SETTING
							--not sh_hsync when others;

--with switch(5 downto 4) select
		out_vsync <= 	--gr_vsync when "00",				-- STABLE SETTING
							--sh_vsync when "01",
							not gr_vsync; -- when "10",
							--not sh_vsync when others;
							
-- 
-- "equivalent" to circuit here: https://cloud.mail.ru/public/FaGH/Jeve8hrKJ/ploca/sch_ttl.png
-- timings reverse engineered from: https://www.futurlec.com/74LS/74LS221.shtml
--h_shot: oneshot Port map ( 
--			trigger => gr_hsync,
--         tick => dotclk,			-- 1 tick is 83.33ns
--         duration => X"00AD", --h_duration, 
--         shot => sh_hsync
--		);
--
--enable_hshot <= '0' when (switch(2 downto 1) = "00") else '0';		
--h_shot_reg: interactivereg Port map ( 
--				reset => RESET,
--				clk => freq2,
--				enable => enable_hshot,
--				init => X"00AD",		-- STABLE SETTING, about 144ms
--				up => button(1),
--				down => button(0),
--				value => open --h_duration
--		);
--
--v_shot: oneshot Port map ( 
--			trigger => gr_vsync,
--         tick => dotclk,			-- 1 tick is 83.33ns
--         duration => X"2000", --v_duration, 	
--         shot => sh_vsync
--		);
--		
--enable_vshot <= '0' when (switch(2 downto 1) = "01") else '0';		
--v_shot_reg: interactivereg Port map ( 
--				reset => RESET,
--				clk => freq2,
--				enable => enable_vshot,
--				init => X"0200", 		-- STABLE SETTING, about 426ms -- NOT USED!
--				up => button(1),
--				down => button(0),
--				value => open --v_duration
--		);
--

leds: fourdigitsevensegled Port map ( 
			-- inputs
			hexdata => hexdata,
			digsel => digsel,
			showdigit => showdigit,
			showdot(3 downto 2) => std_logic_vector(max(9 downto 8)),
			showdot(1 downto 0) => std_logic_vector(min(9 downto 8)),
			-- outputs
			anode => AN,
			segment(7) => DOT,
			segment(6 downto 0) => A_TO_G
		);

showdigit <= "1111"; -- when (data(15) = '1') else (others => freq2); 
----h <= digsel(0) and digsel0_delayed;
--
--cnt_hsync: signalcounter Port map ( 
--				clk => dotclk,
--				reset => RESET,
--				input => out_hsync,
--				sel => switch(0),
--				count => hsync_cnt
--		);
--
--cnt_vsync: signalcounter Port map ( 
--				clk => dotclk,
--				reset => RESET,
--				input => out_vsync,
--				sel => switch(0),
--				count => vsync_cnt
--		);
--

--h_duration <= std_logic_vector(to_unsigned(mouse_x, 16));
--v_duration <= std_logic_vector(to_unsigned(mouse_y, 16));

hexsel <= switch(3 downto 2) & digsel;

with hexsel select
--	hexdata <= 	hsync_cnt(3 downto 0) when "0000",	
--					hsync_cnt(7 downto 4) when "0001",
--					hsync_cnt(11 downto 8) when "0010",
--					hsync_cnt(15 downto 12) when "0011",
--					vsync_cnt(3 downto 0) when "0100",
--					vsync_cnt(7 downto 4) when "0101",
--					vsync_cnt(11 downto 8) when "0110",
--					vsync_cnt(15 downto 12) when "0111",
	hexdata <= 	h_duration(3 downto 0) when "0000",	
					h_duration(7 downto 4) when "0001",
					h_duration(11 downto 8) when "0010",
					h_duration(15 downto 12) when "0011",
					v_duration(3 downto 0) when "0100",
					v_duration(7 downto 4) when "0101",
					v_duration(11 downto 8) when "0110",
					v_duration(15 downto 12) when "0111",
					--
					--data(3 downto 0) when "1000",
					--data(7 downto 4) when "1001",
					--data(11 downto 8) when "1010",
					--data(15 downto 12) when "1011",
					display(3 downto 0) when "1000",
					display(7 downto 4) when "1001",
					display(11 downto 8) when "1010",
					display(15 downto 12) when "1011",
					--DD(3 downto 0) when "1000",
					--DD(7 downto 4) when "1001",
					--D(3 downto 0) when "1010",
					--D(7 downto 4) when "1011",
					A(3 downto 0) when "1100",
					A(7 downto 4) when "1101",
					A(11 downto 8) when "1110",
					A(15 downto 12) when "1111",
					X"0" when others;
					
--testdelay: configurabledelayline Port map (
--				clk => CLK,
--				reset => RESET,
--				init => '1',
--				delay => SW(7 downto 4),
--				signal_in => digsel(0),
--				signal_out => digsel0_delayed
--		);

--
-- UART input coming either directly from USB2UART, or ADC
-- 
--with switch(7 downto 5) select
--		baudrate_x4 <= freq153600 when "111",
--							freq76800 when "110", 
--							freq38400 when "101",
--							freq19200 when "100",		
--							freq9600 when "011",		
--							freq4800 when "010",		
--							freq2400 when "001", 	
--							freq1200 when others;		

with switch(7 downto 5) select
		baudrate_x2 <= freq76800 when "111", 
							freq38400 when "110",
							freq19200 when "101",		
							freq9600 when "100",		
							freq4800 when "011",		
							freq2400 when "010", 	
							freq1200 when "001",
						   freq600 when others;

with switch(7 downto 5) select
		baudrate_x1 <= freq38400 when "111",
							freq19200 when "110",		
							freq9600 when "101",		
							freq4800 when "100",		
							freq2400 when "011", 
							freq1200 when "010",
							freq600  when "001",
							freq300 when others;		
--
--update_cnt: process(audio_level)
--begin
--	if (rising_edge(audio_level)) then
--		adc_count <= std_logic_vector(unsigned(adc_count) + 1);
--	end if;
--end process;
--
--get_rx_analog: process(baudrate_x4, adc_count, adc_old_count)
--begin
--	if (rising_edge(baudrate_x4)) then
--		if (adc_count /= adc_old_count) then
--			rx_analog <= '0'; -- freq x4 detected as at least 1 "zero" crossing happened in t/4 time
--		else
--			rx_analog <= '1';	-- no freq x4 in this t/4 period
--		end if;
--		adc_old_count <= adc_count;
--	end if;
--end process;
--
--rx_digital <= PMOD(6);
--rx <= rx_analog when (switch(1) = '1') else rx_digital;
--
--serin: uart_receiver Port map ( 
--				rx_clk4 => baudrate_x4,
--				reset => RESET,
--				rx => rx,
--				mode => switch(4 downto 2), 
--				frame_active => frame_active,
--				frame_ready => frame_ready, 
--				frame_valid => frame_valid,
--				frame_data => frame_data
--		);
--
--capture_frame: process(RESET, frame_data, frame_ready)
--begin
--	if (RESET = '1') then
--		sr <= X"FFFFFFFF";
--	else
--		if (rising_edge(frame_ready)) then
--			sr <= sr(15 downto 0) & frame_data;
--		end if;
--	end if;
--end process;
--
--AUDIO_OUT_L <= baudrate_x2 when (PMOD(6) = '1') else baudrate_x4;
--AUDIO_OUT_R <= baudrate_x2 when (PMOD(6) = '1') else baudrate_x4;
--	

f_out <= baudrate_x1 when (switch(0) = '0') else baudrate_x2;
AUDIO_OUT_L <= f_out; --baudrate_x2 when (PMOD(6) = '1') else baudrate_x4;
AUDIO_OUT_R <= f_out; --baudrate_x2 when (PMOD(6) = '1') else baudrate_x4;

--f_in_audio <= '0' when (adc_value = X"00") else '1';
f_in <= f_out when (switch(1) = '0') else f_in_audio;

cnt: freqcounter port map (
			reset => RESET,
         clk => freq2,
         freq => f_in,
			bcd => '1',
         value => freq_value
		);
		
display <= std_logic_vector(max(7 downto 0)) & std_logic_vector(min(7 downto 0)) when (switch(1) = '0') else freq_value;
--	sel 	freq	max<<2	min<<2 (diff=1)
--	000	300		C2			28
-- 001	600		C2			28
-- 010	1200		C1			28
-- 011	2400		BF			2C
-- 100	4800		BB			33
-- 101	9600		A8			3B
-- 110	19200		9A			67
-- 111	38400		83			73
-- 1111	76800		80			69
--	sel	freq		max		min (diff=0)	f_out		f_in_audio
--	000	300		49			00					12B		12B
-- 001	600		48			00					257		257
-- 010	1200		48			00					4AE		4AE
-- 011	2400		43			00					95D		0000
-- 100	4800		36			00					12B9		0000
-- 101	9600		03			00					2573		0000
-- 110	19200		03			00					4AE5		0000
-- 111	38400		01			00					95CA		0000
-- 1111	76800		00			00					????		????
--
---------------------------------------------------------------------------------
---- ADC
---------------------------------------------------------------------------------
--  -- Set ADC channel to 0 (audio left) or 1 (audio right)
  adc_channel <= "000"; -- & switch(0);

  adc_clk <= freq24M;
  
  -- Mercury ADC component
  ADC : entity work.MercuryADC
    port map(
      clock    => adc_clk,
      trigger  => adc_trigger,
      diffn    => '0',
      channel  => adc_channel,
      Dout     => adc_dout,
      OutVal   => adc_done,
      adc_miso => ADC_MISO,
      adc_mosi => ADC_MOSI,
      adc_cs   => ADC_CSN,
      adc_clk  => ADC_SCK
      );
--
--  -- ADC sampling process
  sample_adc : process (adc_clk, adc_trigger, adc_dout)
  begin
    if (rising_edge(adc_clk)) then
      -- Sample the ADC continuously
      if (adc_trigger = '1') then  -- Reset the ADC trigger after a single clock cycle
        adc_trigger <= '0';
      else
			if (adc_done = '1') then  -- After a trigger, wait for the ADC's done signal

--				if (adc_dout(9 downto 1) = "000000000") then
--					audio_level <= '0';
--				else
--					audio_level <= '1';
--				end if;
				if (f_in_audio = '0') then
					if (unsigned(adc_dout) /= "0000000000") then
						f_in_audio <= '1';
					end if;
				else
					if (adc_dout = "0000000000") then
						f_in_audio <= '0';
					end if;
				end if;
				adc_value <= adc_dout(9 downto 2);
					
				if (unsigned(adc_dout) > max) then
					max <= unsigned(adc_dout);
				end if;

				if (unsigned(adc_dout) < min) then
					min <= unsigned(adc_dout);
				end if;

				adc_trigger  <= '1';            -- Request another sample
			end if;
		end if;
    end if;
  end process;

--display <= sr(15 downto 0) when (switch(0) = '0') else freq_value;
--debug <= std_logic_vector(max(9 downto 2)) & std_logic_vector(min(9 downto 2)) when (switch(0) = '0') else freq_value;

end;
