----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:01:38 03/01/2021 
-- Design Name: 
-- Module Name:    vdp_sampler2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity vdp_sampler2 is
    Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           hsync : in  STD_LOGIC;
           vsync : in  STD_LOGIC;
			  pixclk: in STD_LOGIC;
           r : in  STD_LOGIC;
           g : in  STD_LOGIC;
			  b : in  STD_LOGIC;
           a : out  STD_LOGIC_VECTOR (14 downto 0);
           d : out  STD_LOGIC_VECTOR (7 downto 0);
			  limit: in STD_LOGIC_VECTOR (5 downto 0);
			  we_in: in STD_LOGIC;
           we_out : out  STD_LOGIC);
end vdp_sampler2;

architecture Behavioral of vdp_sampler2 is


signal h, h_off: std_logic_vector(8 downto 0);
signal v, v_off: std_logic_vector(8 downto 0);
signal sample: std_logic_vector(7 downto 0);
signal h_ok, v_ok, write_clk: std_logic;
signal cnt, sample_cnt, write_cnt: integer range 0 to 63;

begin

-- output signals
d <= sample;
a <= v_off(7 downto 0) & h_off(7 downto 1);
we_out <= h(0) and write_clk and (not hsync) and (not h_off(8)) and (not v_off(8));

-- offset to ignore all before real pixel data comes in
h_off <= std_logic_vector(unsigned(h) - 27);
v_off <= std_logic_vector(unsigned(v) - 27);
v_ok <= '0' when (unsigned(v_off) > 191) else '1';

-- when to take the sample within the pixel clock period
sample_cnt 	<= to_integer(unsigned(limit(5 downto 0)));
write_cnt 	<= sample_cnt + 2;

-- generate single write pulse
write_clk <= '1' when (write_cnt = cnt) else '0';

on_clk: process(clk, pixclk, cnt, r, g, b)
begin 
	if (pixclk = '0') then
		cnt <= 0;
	else
		if (rising_edge(clk)) then
			cnt <= cnt + 1;
			if (cnt = sample_cnt) then
				sample <= sample(3 downto 0) & '0' & r & g & b;
			end if;
		end if;
	end if;
end process;

on_write_clk: process(write_clk, reset, hsync, h)
begin
	if ((reset or hsync) = '1') then
		h <= "000000000";
	else
		if (rising_edge(write_clk)) then
			h <= std_logic_vector(unsigned(h) + 1);
		end if;
	end if;
end process;

on_hsync: process(hsync, reset, vsync, v)
begin
	if ((reset or vsync) = '1') then
		v <= "000000000";
	else
		if (falling_edge(hsync)) then
			v <= std_logic_vector(unsigned(v) + 1);
		end if;
	end if;
end process;

end Behavioral;

