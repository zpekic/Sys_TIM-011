----------------------------------------------------------------------------------
-- Company: @Home
-- Engineer: zpekic@hotmail.com
-- 
-- Create Date: 08/29/2020 11:13:02 PM
-- Design Name: Various TIM-011 components
-- Module Name: sys_tim-011_mercury - Behavioral
-- Project Name: 
-- Target Devices: https://www.micro-nova.com/mercury/ + Baseboard
-- Input devices: 
--
-- Tool Versions: ISE 14.7 (nt)
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.99 - Kinda works...
-- Additional Comments:
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
--use work.tms0800_package.all;

entity sys_tim011_mercury is
    Port ( 
				-- 50MHz on the Mercury board
				CLK: in std_logic;
				
				-- 12MHz external clock
				EXT_CLK: in std_logic;
				
				-- Master reset button on Mercury board
				USR_BTN: in std_logic; 

				-- Switches on baseboard
				-- SW(0) -- direction when scrolling
				-- SW(1) -- data source selection for 7seg display
				-- SW(2) -- palette selection (best on)
				-- SW(3) -- palette selection (best off)
				-- SW(4) -- off
				-- SW(5) -- on
				-- SW(6) -- off
				-- SW(7)	-- off

				SW: in std_logic_vector(7 downto 0); 

				-- Push buttons on baseboard
				-- BTN0 - scroll
				-- BTN1 - video only test pattern (memory not affected)
				-- BTN2 - fill left/right
				-- BTN3 - fill top/down
				BTN: in std_logic_vector(3 downto 0); 

				-- Stereo audio output on baseboard
				--AUDIO_OUT_L, AUDIO_OUT_R: out std_logic;

				-- 7seg LED on baseboard 
				A_TO_G: out std_logic_vector(6 downto 0); 
				AN: out std_logic_vector(3 downto 0); 
				DOT: out std_logic; 
				-- 4 LEDs on Mercury board (3 and 2 are used by VGA VSYNC and HSYNC)
				--LED: inout std_logic_vector(3 downto 0);

				-- ADC interface
				-- channel	input
				-- 0			Audio Left
				-- 1 			Audio Right
				-- 2			Temperature
				-- 3			Light	
				-- 4			Pot
				-- 5			Channel 5 (free)
				-- 6			Channel 6 (free)
				-- 7			Channel 7 (free)
				--ADC_MISO: in std_logic;
				--ADC_MOSI: out std_logic;
				--ADC_SCK: out std_logic;
				--ADC_CSN: out std_logic;
				PS2_DATA: inout std_logic;
				PS2_CLOCK: inout std_logic;

				--VGA interface
				--register state is traced to VGA after each instruction if SW0 = on
				--640*480 50Hz mode is used, which give 80*60 character display
				--but to save memory, only 80*50 are used which fits into 4k video RAM
				HSYNC: out std_logic;
				VSYNC: out std_logic;
				RED: out std_logic_vector(2 downto 0);
				GRN: out std_logic_vector(2 downto 0);
				BLU: out std_logic_vector(1 downto 0);
				
				--PMOD interface
				--connection to https://store.digilentinc.com/pmod-kypd-16-button-keypad/
				PMOD: inout std_logic_vector(7 downto 0)
          );
end sys_tim011_mercury;

architecture Structural of sys_tim011_mercury is

component Grafika is
    Port ( -- 
	 		  dotclk : in  STD_LOGIC;
           a : in  STD_LOGIC_VECTOR (15 downto 0);
           nRD : in  STD_LOGIC;
           nWR : in  STD_LOGIC;
           d : inout  STD_LOGIC_VECTOR (7 downto 0);
           ioe : in  STD_LOGIC;
           nScroll : in  STD_LOGIC;
			  -- debug
			  test: in STD_LOGIC;
			  vid_gated: STD_LOGIC;
			  -- monitor side
			  hsync: out STD_LOGIC;
			  vsync: out STD_LOGIC;
			  vid1: out STD_LOGIC;
			  vid2: out STD_LOGIC
			);
end component;

component oneshot is
    Port ( trigger : in  STD_LOGIC;
           tick : in  STD_LOGIC;
           duration : in  STD_LOGIC_VECTOR (15 downto 0);
           shot : out  STD_LOGIC);
end component;

component sn74ls283 is
    Port ( c0 : in  STD_LOGIC;
           a : in  STD_LOGIC_VECTOR (4 downto 1);
           b : in  STD_LOGIC_VECTOR (4 downto 1);
           s : out  STD_LOGIC_VECTOR (4 downto 1);
           c4 : out  STD_LOGIC);
end component;

component sn74ls374 is
    Port ( nOC : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           D : in  STD_LOGIC_VECTOR (7 downto 0);
           Q : out  STD_LOGIC_VECTOR (7 downto 0));
end component;

component sn74hc4040 is
    Port ( q12_1 : out  STD_LOGIC;
           q6_2 : out  STD_LOGIC;
           q5_3 : out  STD_LOGIC;
           q7_4 : out  STD_LOGIC;
           q4_5 : out  STD_LOGIC;
           q3_6 : out  STD_LOGIC;
           q2_7 : out  STD_LOGIC;
           q1_9 : out  STD_LOGIC;
           clock_10 : in  STD_LOGIC;
           reset_11 : in  STD_LOGIC;
           q9_12 : out  STD_LOGIC;
           q8_13 : out  STD_LOGIC;
           q10_14 : out  STD_LOGIC;
           q11_15 : out  STD_LOGIC);
end component;

component fourdigitsevensegled is
    Port ( -- inputs
			  hexdata : in  STD_LOGIC_VECTOR (3 downto 0);
           digsel : in  STD_LOGIC_VECTOR (1 downto 0);
           showdigit : in  STD_LOGIC_VECTOR (3 downto 0);
           showdot : in  STD_LOGIC_VECTOR (3 downto 0);
			  -- outputs
           anode : out  STD_LOGIC_VECTOR (3 downto 0);
           segment : out  STD_LOGIC_VECTOR (7 downto 0)
			 );
end component;

component interactivereg is
    Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           enable : in  STD_LOGIC;
           init : in  STD_LOGIC_VECTOR (15 downto 0);
           up : in  STD_LOGIC;
           down : in  STD_LOGIC;
           value : buffer  STD_LOGIC_VECTOR (15 downto 0));
end component;

component freqcounter is
    Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           freq : in  STD_LOGIC;
			  bcd:	in STD_LOGIC;
			  double: in STD_LOGIC;
			  limit: in STD_LOGIC_VECTOR(15 downto 0);
			  ge: out STD_LOGIC;
           value : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component uart_receiver is
    Port ( rx_clk4 : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           rx : in  STD_LOGIC;
           mode : in  STD_LOGIC_VECTOR (2 downto 0);
			  frame_active: out  STD_LOGIC;
           frame_ready : out  STD_LOGIC;
           frame_valid : out  STD_LOGIC;
           frame_data : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component uart_sender is
	 Port (  tx_clk  : in  STD_LOGIC;
				reset  : in  STD_LOGIC;
				tx  : out  STD_LOGIC;
				ready: out STD_LOGIC;
				mode : in  STD_LOGIC_VECTOR (2 downto 0); 
				send : in  STD_LOGIC; 
				enable : in  STD_LOGIC;
				data : in STD_LOGIC_VECTOR(7 downto 0));
end component;
		
component signalcounter is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           input : in  STD_LOGIC;
           sel : in  STD_LOGIC;
           count : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component configurabledelayline is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           init : in  STD_LOGIC;
           delay : in  STD_LOGIC_VECTOR (3 downto 0);
           signal_in : in  STD_LOGIC;
           signal_out : out  STD_LOGIC);
end component;

component vga_controller is
    Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           hsync : out  STD_LOGIC;
           vsync : out  STD_LOGIC;
			  x_valid: out STD_LOGIC;
			  y_valid: out STD_LOGIC;
			  h_active: out STD_LOGIC;
			  v_active: out STD_LOGIC;
           x : out  STD_LOGIC_VECTOR (8 downto 0);
           y : out  STD_LOGIC_VECTOR (7 downto 0));
end component;

--component rx_reg is
--    Port ( clk : in  STD_LOGIC;
--           reset : in  STD_LOGIC;
--           enable : in  STD_LOGIC;
--           rx : in  STD_LOGIC;
--           d : out  STD_LOGIC_VECTOR (7 downto 0);
--           dready : out  STD_LOGIC);
--end component;

--component tapeuart is
--    Port ( reset : in  STD_LOGIC;
--           serout : out  STD_LOGIC;
--           serin : in  STD_LOGIC;
--			  freq_mark: in STD_LOGIC;
--			  freq_space: in STD_LOGIC;
--           audio_left : out  STD_LOGIC;
--           audio_right : out  STD_LOGIC;
--           adc_clk : in  STD_LOGIC;
--           adc_samplefreq : in  STD_LOGIC;
--           adc_miso : in  STD_LOGIC;
--           adc_mosi : out  STD_LOGIC;
--           adc_sck : out  STD_LOGIC;
--           adc_csn : out  STD_LOGIC;
--			  --
--			  debugsel: in STD_LOGIC;
--			  debug: out STD_LOGIC_VECTOR(15 downto 0)
--			);
--end component;

--component memconsole is
--    Port ( clk : in  STD_LOGIC;
--           reset : in  STD_LOGIC;
--           control : in  STD_LOGIC_VECTOR (3 downto 0);
--           EN : out  STD_LOGIC;
--           RD : out  STD_LOGIC;
--           WR : out  STD_LOGIC;
--           A : out  STD_LOGIC_VECTOR (15 downto 0);
--           D : inout  STD_LOGIC_VECTOR (7 downto 0);
--           DD : out  STD_LOGIC_VECTOR (7 downto 0));
--end component;

component ps2tim is
    Port ( reset : in  STD_LOGIC;
           uart_clk4 : in  STD_LOGIC;
           uart_rx : in  STD_LOGIC;
           uart_tx : out  STD_LOGIC;
			  uart_mode: in STD_LOGIC_VECTOR(2 downto 0);
           ps2_clk : inout  STD_LOGIC;
           ps2_data : inout  STD_LOGIC;
			  kbd_alt: buffer STD_LOGIC;
			  kbd_shift: buffer STD_LOGIC;
			  kbd_ctrl: buffer STD_LOGIC;
			  kbd_caps: buffer STD_LOGIC;
			  debugsel: in STD_LOGIC;
           debug : out  STD_LOGIC_VECTOR (15 downto 0));
end component;

component debouncer8channel is
    Port ( clock : in STD_LOGIC;
           reset : in STD_LOGIC;
           signal_raw : in STD_LOGIC_VECTOR (7 downto 0);
           signal_debounced : out STD_LOGIC_VECTOR (7 downto 0));
end component;



component ram32k8 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END component;

--component memtester is
--    Port ( clk : in  STD_LOGIC;
--           reset : in  STD_LOGIC;
--			  fill: in STD_LOGIC;
--			  direction: in STD_LOGIC;
--           EN : out  STD_LOGIC;
--           RD : out  STD_LOGIC;
--           WR : out  STD_LOGIC;
--           A : out  STD_LOGIC_VECTOR (15 downto 0);
--           D : inout  STD_LOGIC_VECTOR (7 downto 0);
--           DD : out  STD_LOGIC_VECTOR (7 downto 0));
--end component;
--
--type palette is array (0 to 15) of std_logic_vector(2 downto 0);
--signal bgr: palette := (
--	"011",	-- yellow -- this palette looks bad probably because base background color is not black
--	"110",	-- cyan
--	"101",	-- purple
--	"111",	-- white
--
--	"000",	-- black
--	"101",	-- purple
--	"110",	-- cyan
--	"100",	-- blue
--
--	"000",	-- black
--	"011",	-- yellow
--	"110",	-- cyan
--	"010",	-- green
--
--	"000",	-- black
--	"011",	-- yellow
--	"101",	-- purple
--	"001" 	-- red
--);

type vga_palette is array (0 to 15) of std_logic_vector(7 downto 0);
signal rgb: vga_palette := (
	"00000011", -- screen outside of TIM window
	"00000011", -- screen outside of TIM window
	"00000011", -- screen outside of TIM window
	"00000011", -- screen outside of TIM window
	"00011100", -- screen outside of TIM window
	"00011100", -- screen outside of TIM window
	"00011100", -- screen outside of TIM window
	"00011100", -- screen outside of TIM window
	"11100000", -- screen outside of TIM window
	"11100000", -- screen outside of TIM window
	"11100000", -- screen outside of TIM window
	"11100000", -- screen outside of TIM window
	"00000000", -- black
	"01001001", -- dk gray
	"10010010", -- lt gray
	"11111111"  -- white
);

signal RESET: std_logic;

-- debug
signal digsel: std_logic_vector(1 downto 0);
signal hexdata, hexsel, showdigit: std_logic_vector(3 downto 0);
---

--- frequency signals
signal freq24M, freq25M, dotclk, freq0M75: std_logic;
signal prescale_baud, prescale_power: integer range 0 to 65535;
signal freq153600, freq76800, freq38400, freq19200, freq9600, freq4800, freq2400, freq1200, freq600, freq300, freq150: std_logic;		
signal freq4096, freq2, freq4: std_logic;		

--- video sync signals
signal x_valid, y_valid: std_logic;
signal h_active, v_active : std_logic;
signal vga_x: std_logic_vector(8 downto 0); -- 512 pixels horizontally
signal vga_y: std_logic_vector(7 downto 0); -- 256 pixels vertically
-- video data signals
signal color_index: std_logic_vector(3 downto 0);
signal vga_color: std_logic_vector(7 downto 0);
signal pair: std_logic_vector(1 downto 0); -- 2 bit pixel
-- video memory bus
signal vram_wr_nrd, tim_wr_nrd: std_logic;
signal vram_dina, vram_douta: std_logic_vector(7 downto 0);
signal vram_addra, vga_a, tim_a: std_logic_vector(14 downto 0);
signal vram_wea: std_logic_vector(0 downto 0);

---
signal switch, button: std_logic_vector(7 downto 0);


--alias ps2_data: std_logic is LED(0);
--alias ps2_clk: std_logic is LED(1);

-- UART
signal frame_ready, frame_valid, frame_active: std_logic;
signal frame_data, uart_frame, display: std_logic_vector(15 downto 0);
--signal rx, rx_analog, rx_digital: std_logic;
signal baudrate_x1, baudrate_x2, baudrate_x4: std_logic;
signal sr: std_logic_vector(31 downto 0);

signal kbd_alt, kbd_shift, kbd_ctrl, kbd_caps: STD_LOGIC;

-- https://reference.digilentinc.com/reference/pmod/pmodusbuart/reference-manual
alias nRTS: std_logic is PMOD(4); 	-- out, active low
alias RXD_TTY: std_logic is PMOD(5);		-- in
alias TXD_TTY: std_logic is PMOD(6);		-- out
alias nCTS: std_logic is PMOD(7);	-- in, active low

begin
   
-- connect to "oscilloscope"
PMOD(0) <= baudrate_x4;
PMOD(1) <= baudrate_x1;
PMOD(2) <= RXD_TTY;
PMOD(3) <= TXD_TTY;
	
RESET <= USR_BTN;
	
clockgen: sn74hc4040 port map (
			clock_10 => EXT_CLK,	-- 48MHz "half-size" crystal on Mercury baseboard
			reset_11 => RESET,
			q1_9 => freq24M, 
			q2_7 => dotclk,
			q3_6 => open, --PMOD(7),			-- 6
			q4_5 => open, --PMOD(6),			-- 3
			q5_3 => open, --PMOD(5),			-- 1.5
			q6_2 => freq0M75, --PMOD(4), 		-- 0.75
			q7_4 =>   open,		-- 0.325
			q8_13 =>  open,		-- 0.1625
			q9_12 =>  open,		-- 0.08125
			q10_14 => open,		-- 0.040625
			q11_15 => digsel(0),	-- 0.0203125
			q12_1 =>  digsel(1)	-- 0.01015625
		);
--
prescale: process(CLK, freq153600, freq4096)
begin
	if (rising_edge(CLK)) then
		freq25M <= not freq25M;	-- used for VGA 640*480
		if (prescale_baud = 0) then
			freq153600 <= not freq153600;
			prescale_baud <= (50000000 / (2 * 153600));
		else
			prescale_baud <= prescale_baud - 1;
		end if;
		if (prescale_power = 0) then
			freq4096 <= not freq4096;
			prescale_power <= (50000000 / (2 * 4096));
		else
			prescale_power <= prescale_power - 1;
		end if;
	end if;
end process;
--
baudgen: sn74hc4040 port map (
			clock_10 => freq153600,
			reset_11 => RESET,
			q1_9 => freq76800, 
			q2_7 => freq38400,
			q3_6 => freq19200,		
			q4_5 => freq9600,		
			q5_3 => freq4800,		
			q6_2 => freq2400, 	
			q7_4 => freq1200,		
			q8_13 => freq600,		
			q9_12 =>  freq300,
			q10_14 => freq150,	
			q11_15 => open,	
			q12_1 =>  open	
		);
--
powergen: sn74hc4040 port map (
			clock_10 => freq4096,
			reset_11 => RESET,
			q1_9 => open, 
			q2_7 => open,
			q3_6 => open,		
			q4_5 => open,		
			q5_3 => open,		
			q6_2 => open, 	
			q7_4 => open,		
			q8_13 => open,		
			q9_12 =>  open,	
			q10_14 => freq4,	
			q11_15 => freq2,	
			q12_1 =>  open	
		);
--	
	debounce_sw: debouncer8channel Port map ( 
		clock => freq19200, 
		reset => RESET,
		signal_raw => SW,
		signal_debounced => switch
	);

	debounce_btn: debouncer8channel Port map ( 
		clock => freq19200, 
		reset => RESET,
		signal_raw(7 downto 4) => "0000",
		signal_raw(3 downto 0) => BTN,
		signal_debounced => button
	);
	
kbd: ps2tim Port map ( 
			reset => RESET,
         uart_clk4 => baudrate_x4, -- baudrate = /4 = 9600
         uart_rx => TXD_TTY,
         uart_tx => RXD_TTY,
			uart_mode => switch(4 downto 2),
         ps2_clk => PS2_CLOCK, --LED(1),
         ps2_data => PS2_DATA, --LED(0),
			kbd_alt => kbd_alt,
			kbd_shift => kbd_shift,
			kbd_ctrl => kbd_ctrl,
			kbd_caps => kbd_caps,
			debugsel => switch(0),
         debug => display
		);

vga: vga_controller Port map ( 
		reset => RESET,
      clk => freq25M,
      hsync => HSYNC,
      vsync => VSYNC,
		x_valid => x_valid,
		y_valid => y_valid,
		h_active => open,
		v_active => open,
      x => vga_x,
      y => vga_y
	);

mem: ram32k8 PORT MAP (
    clka => CLK,
	 ena => '1',
    wea => vram_wea,
    addra => vram_addra,
    dina => vram_dina,
    douta => vram_douta
  );

vram_wr_nrd <= '0'; --'0' when (y_valid = '1') else tim_rd_nwr;

vram_addra <= (vga_y & vga_x(8 downto 2)) when (y_valid = '1') else tim_a;
vram_wea <= (others => vram_wr_nrd);

-- pixels are stored 11003322
-- see https://github.com/zpekic/Sys_TIM-011/blob/master/Img2Tim/Img2Tim/Program.cs
with vga_x(1 downto 0) select pair <=
	vram_douta(5 downto 4) when "00",
	vram_douta(7 downto 6) when "01",
	vram_douta(1 downto 0) when "10",
	vram_douta(3 downto 2) when others;

-- color index also takes into account selected palette and if in TIM window
color_index <= y_valid & x_valid & pair; 

-- now convert to VGA 8-bit color
vga_color <= rgb(to_integer(unsigned(color_index)));
RED <= vga_color(7 downto 5);
GRN <= vga_color(4 downto 2);
BLU <= vga_color(1 downto 0);

--console: memconsole Port map(
--			clk => freq2,
--         reset => RESET,
--         control => button(3 downto 0),
--         EN => vm_en,
--         RD => vm_rd,
--         WR => vm_wr,
--         A => A,
--         D => D,
--         DD => DD
--	);

--mtest: memtester Port map(
--			clk => test_clk,
--         reset => RESET,
--			fill => test_dynamic,
--			direction => button(2),
--         EN => vm_en,
--         RD => vm_rd,
--         WR => vm_wr,
--         A => A,
--         D => D,
--         DD => DD
--	);
----	
--test_static <= '1' when (button(3 downto 0) = "0010") else '0';
--test_dynamic <= '0' when (button(3 downto 2) = "00") else '1';
--test_scroll <= nScrollEnable when (button(3 downto 0) = "0001") else '1';
--
--test_clk <= freq38400 when (button(3 downto 2) = "11") else freq9600;
--
---- scroll logic
--nScrollEnable <= vm_en or vm_rd or vm_wr;	-- low if all all, meaning no other bus activity
--
--offset_reg: sn74ls374 Port map ( 
--			nOC => nScrollEnable,
--         CLK => test_scroll,
--         D => offset_new,
--         Q => D
--	);
--
--offset_add_hi: sn74ls283 Port map ( -- add +1 or -1 to offset)
--			c0 => offset_add_lo_cout,
--			a(4) => switch(0),
--			a(3) => switch(0),
--			a(2) => switch(0),
--			a(1) => switch(0),
--			b => D(7 downto 4),
--			s => offset_new(7 downto 4),
--			c4 => open
--	);
--	
--offset_add_lo: sn74ls283 Port map ( 
--			c0 => '0',
--			a(4) => switch(0),
--			a(3) => switch(0),
--			a(2) => switch(0),
--			a(1) => '1',
--			b => D(3 downto 0),
--			s => offset_new(3 downto 0),
--			c4 => offset_add_lo_cout
--	);	
--	

--	video: Grafika port map (
--		-- system
--		  dotclk => dotclk,
--		  A(15) => '1',	-- mapped to 0x8000 - 0xFFFF or extended IO space
--		  A(14 downto 0) => A(14 downto 0),
--		  nRD => not (vm_rd),
--		  nWR => not (vm_wr),
--		  d => D,
--		  ioe => vm_en,
--		  nScroll => test_scroll,
--		-- debug
--		  test => test_static,
--		  vid_gated => '0', -- do not gate vid1/2 on dotclk (this is different from original!)
--		-- monitor side
--		  hsync => gr_hsync, --HSYNC,
--		  vsync => gr_vsync,--VSYNC,
--		  vid1 => gr_vid1, --BLU(0),
--		  vid2 => gr_vid2  --BLU(1)
--	);
	
--LED(0) <= dotclk;
--LED(1) <= vm_en;
--LED(2) <= x_valid;
--LED(3) <= y_valid;

-- Connect to GBS8200 gray wire
	--PMOD(3) <= out_hsync xor out_vsync;
	
-- connect to GBS8200 blue / green / red wires
	--PMOD(2 downto 0) <= bgr(to_integer(unsigned(color)));
	--color <= switch(3 downto 2) & gr_vid2 & gr_vid1;

--	HSYNC <= not sh_hsync;
--	VSYNC <= not sh_vsync;
--	BLU(1) <= switch(1) xor gr_vid2;
--	BLU(0) <= switch(0) xor gr_vid1;
--	RED <= "000";
--	GRN <= "000";

--with switch(7 downto 6) select
		--out_hsync <= 	gr_hsync; -- when "00",
							--sh_hsync when "01",
							--not gr_hsync when "10",			-- STABLE SETTING
							--not sh_hsync when others;

--with switch(5 downto 4) select
		--out_vsync <= 	--gr_vsync when "00",				-- STABLE SETTING
							--sh_vsync when "01",
							--not gr_vsync; -- when "10",
							--not sh_vsync when others;
							
leds: fourdigitsevensegled Port map ( 
			-- inputs
			hexdata => hexdata,
			digsel => digsel,
			showdigit => showdigit,
			--showdot(3) => "00", --std_logic_vector(max(9 downto 8)),
			--showdot(2) => "00", --std_logic_vector(min(9 downto 8)),
			showdot(3) => kbd_alt,
			showdot(2) => kbd_shift,
			showdot(1) => kbd_ctrl,
			showdot(0) => kbd_caps,
			-- outputs
			anode => AN,
			segment(7) => DOT,
			segment(6 downto 0) => A_TO_G
		);

showdigit <= "1111"; -- when (data(15) = '1') else (others => freq2); 

with digsel select
	hexdata <= 	display(3 downto 0) when "00",	
					display(7 downto 4) when "01",
					display(11 downto 8) when "10",
					display(15 downto 12) when others;

--
-- UART input coming either directly from USB2UART, or ADC
-- 
with switch(7 downto 5) select
		baudrate_x4 <= freq153600 when "111",
							freq76800 when "110", 
							freq38400 when "101",
							freq19200 when "100",		
							freq9600 when "011",		
							freq4800 when "010",		
							freq2400 when "001", 	
							freq1200 when others;		

with switch(7 downto 5) select
		baudrate_x2 <= freq76800 when "111", 
							freq38400 when "110",
							freq19200 when "101",		
							freq9600 when "100",		
							freq4800 when "011",		
							freq2400 when "010", 	
							freq1200 when "001",
						   freq600 when others;

with switch(7 downto 5) select
		baudrate_x1 <= freq38400 when "111",
							freq19200 when "110",		
							freq9600 when "101",		
							freq4800 when "100",		
							freq2400 when "011", 
							freq1200 when "010",
							freq600  when "001",
							freq300 when others;		

--streamer: tapeuart port map ( 
--				reset => RESET,
--				serout => open, --RXD_TTY,
--				serin => '1', --TXD_TTY,
--				freq_mark => freq4800,
--				freq_space => freq2400,
--				audio_left => AUDIO_OUT_L,
--				audio_right => AUDIO_OUT_R,
--				adc_clk => freq24M,
--				adc_samplefreq => freq0M75,
--				adc_miso => ADC_MISO,
--				adc_mosi => ADC_MOSI,
--				adc_sck => ADC_SCK,
--				adc_csn => ADC_CSN,
--				----
--				debugsel => switch(0),
--				debug => open --display
--			);

--
--serin: uart_receiver Port map ( 
--				rx_clk4 => baudrate_x4,
--				reset => RESET,
--				rx => RXD_TTY,	-- "txd" looking from the sender side
--				mode => switch(4 downto 2), 
--				frame_active => frame_active,
--				frame_ready => frame_ready, 
--				frame_valid => frame_valid,
--				frame_data => frame_data
--		);
--
--capture_frame: process(RESET, frame_data, frame_ready)
--begin
--	if (RESET = '1') then
--		sr <= X"FFFFFFFF";
--	else
--		if (rising_edge(frame_ready)) then
--			sr <= sr(15 downto 0) & frame_data;
--		end if;
--	end if;
--end process;

--serout: uart_sender port map (
--				tx_clk => baudrate_x1,
--				reset => RESET,
--				tx => RXD_TTY,	-- "rxd" looking from the receiver side
--				ready => open,
--				mode => switch(4 downto 2), 
--				send => frame_ready, 
--				enable => frame_valid,
--				data => frame_data(7 downto 0)
--		);

----display <= std_logic_vector(max(7 downto 0)) & std_logic_vector(min(7 downto 0)) when (switch(1) = '0') else freq_value;
--display <= freq_value;
--	sel 	freq	max<<2	min<<2 (diff=1)
--	000	300		C2			28
-- 001	600		C2			28
-- 010	1200		C1			28
-- 011	2400		BF			2C
-- 100	4800		BB			33
-- 101	9600		A8			3B
-- 110	19200		9A			67
-- 111	38400		83			73
-- 1111	76800		80			69
--	sel	freq		max		min (diff=0)	f_out		f_in_audio
--	000	300		49			00					12B		12B
-- 001	600		48			00					257		257
-- 010	1200		48			00					4AE		4AE
-- 011	2400		43			00					95D		0000
-- 100	4800		36			00					12B9		0000
-- 101	9600		03			00					2573		0000
-- 110	19200		03			00					4AE5		0000
-- 111	38400		01			00					95CA		0000
-- 1111	76800		00			00					????		????
--
		
--
--  -- ADC sampling process
--  sample_adc : process (adc_clk, adc_trigger, adc_dout)
--  begin
--    if (rising_edge(adc_clk)) then
--      -- Sample the ADC continuously
--      if (adc_trigger = '1') then  -- Reset the ADC trigger after a single clock cycle
--        adc_trigger <= '0';
--      end if;
--		
--		if (adc_done = '1') then  -- After a trigger, wait for the ADC's done signal
--
----				if (adc_dout(9 downto 1) = "000000000") then
----					audio_level <= '0';
----				else
----					audio_level <= '1';
----				end if;
--			if (f_in_audio = '0') then
--				if (unsigned(adc_dout) > "0000100100") then
--					f_in_audio <= '1';
--				end if;
--			else
--				if (unsigned(adc_dout) < "0000100100") then
--					f_in_audio <= '0';
--				end if;
--			end if;
--			adc_value <= adc_dout(9 downto 2);
--				
--			if (unsigned(adc_dout) > max) then
--				max <= unsigned(adc_dout);
--			end if;
--
--			if (unsigned(adc_dout) < min) then
--				min <= unsigned(adc_dout);
--			end if;
--
--			adc_trigger  <= '1';            -- Request another sample
--		end if;
--    end if;
--  end process;

--hexsel <= switch(3 downto 2) & digsel;
--
--with hexsel select
----	hexdata <= 	hsync_cnt(3 downto 0) when "0000",	
----					hsync_cnt(7 downto 4) when "0001",
----					hsync_cnt(11 downto 8) when "0010",
----					hsync_cnt(15 downto 12) when "0011",
----					vsync_cnt(3 downto 0) when "0100",
----					vsync_cnt(7 downto 4) when "0101",
----					vsync_cnt(11 downto 8) when "0110",
----					vsync_cnt(15 downto 12) when "0111",
--	hexdata <= 	h_duration(3 downto 0) when "0000",	
--					h_duration(7 downto 4) when "0001",
--					h_duration(11 downto 8) when "0010",
--					h_duration(15 downto 12) when "0011",
--					v_duration(3 downto 0) when "0100",
--					v_duration(7 downto 4) when "0101",
--					v_duration(11 downto 8) when "0110",
--					v_duration(15 downto 12) when "0111",
--					--
--					--data(3 downto 0) when "1000",
--					--data(7 downto 4) when "1001",
--					--data(11 downto 8) when "1010",
--					--data(15 downto 12) when "1011",
--					display(3 downto 0) when "1000",
--					display(7 downto 4) when "1001",
--					display(11 downto 8) when "1010",
--					display(15 downto 12) when "1011",
--					--DD(3 downto 0) when "1000",
--					--DD(7 downto 4) when "1001",
--					--D(3 downto 0) when "1010",
--					--D(7 downto 4) when "1011",
--					std_logic_vector(min(3 downto 0)) when "1100",
--					std_logic_vector(min(7 downto 4)) when "1101",
--					std_logic_vector(max(3 downto 0)) when "1110",
--					std_logic_vector(max(7 downto 4)) when "1111",
--					X"0" when others;

--display <= freq_value; --sr(15 downto 0);

--display <= sr(15 downto 0) when (switch(0) = '0') else freq_value;
--debug <= std_logic_vector(max(9 downto 2)) & std_logic_vector(min(9 downto 2)) when (switch(0) = '0') else freq_value;

----h <= digsel(0) and digsel0_delayed;
--
--cnt_hsync: signalcounter Port map ( 
--				clk => dotclk,
--				reset => RESET,
--				input => out_hsync,
--				sel => switch(0),
--				count => hsync_cnt
--		);
--
--cnt_vsync: signalcounter Port map ( 
--				clk => dotclk,
--				reset => RESET,
--				input => out_vsync,
--				sel => switch(0),
--				count => vsync_cnt
--		);
--

--h_duration <= std_logic_vector(to_unsigned(mouse_x, 16));
--v_duration <= std_logic_vector(to_unsigned(mouse_y, 16));

-- 
-- "equivalent" to circuit here: https://cloud.mail.ru/public/FaGH/Jeve8hrKJ/ploca/sch_ttl.png
-- timings reverse engineered from: https://www.futurlec.com/74LS/74LS221.shtml
--h_shot: oneshot Port map ( 
--			trigger => gr_hsync,
--         tick => dotclk,			-- 1 tick is 83.33ns
--         duration => X"00AD", --h_duration, 
--         shot => sh_hsync
--		);
--
--enable_hshot <= '0' when (switch(2 downto 1) = "00") else '0';		
--h_shot_reg: interactivereg Port map ( 
--				reset => RESET,
--				clk => freq2,
--				enable => enable_hshot,
--				init => X"00AD",		-- STABLE SETTING, about 144ms
--				up => button(1),
--				down => button(0),
--				value => open --h_duration
--		);
--
--v_shot: oneshot Port map ( 
--			trigger => gr_vsync,
--         tick => dotclk,			-- 1 tick is 83.33ns
--         duration => X"2000", --v_duration, 	
--         shot => sh_vsync
--		);
--		
--enable_vshot <= '0' when (switch(2 downto 1) = "01") else '0';		
--v_shot_reg: interactivereg Port map ( 
--				reset => RESET,
--				clk => freq2,
--				enable => enable_vshot,
--				init => X"0200", 		-- STABLE SETTING, about 426ms -- NOT USED!
--				up => button(1),
--				down => button(0),
--				value => open --v_duration
--		);
--

--testdelay: configurabledelayline Port map (
--				clk => CLK,
--				reset => RESET,
--				init => '1',
--				delay => SW(7 downto 4),
--				signal_in => digsel(0),
--				signal_out => digsel0_delayed
--		);

end;
